module 4xSA_Cache(
    input clk,
    input rst,
);
